module top_module(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);
    wire carry1, carry2;
    add16 low_16(a[15:0], b[15:0], 1'b0, sum[15:0], carry1);
    add16 high_16(a[31:16], b[31:16], carry1, sum[31:16], carry2);
endmodule